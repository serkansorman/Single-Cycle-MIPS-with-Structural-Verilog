module addop(sum,x,y,cout);
input [31:0] x,y;
output cout;
output[31:0] sum;
wire ov,c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29,c30,c31;

full_adder fa1(x[0],y[0],1'b0,sum[0],c1);
full_adder fa2(x[1],y[1],c1,sum[1],c2);
full_adder fa3(x[2],y[2],c2,sum[2],c3);
full_adder fa4(x[3],y[3],c3,sum[3],c4);
full_adder fa5(x[4],y[4],c4,sum[4],c5);
full_adder fa6(x[5],y[5],c5,sum[5],c6);
full_adder fa7(x[6],y[6],c6,sum[6],c7);
full_adder fa8(x[7],y[7],c7,sum[7],c8);
full_adder fa9(x[8],y[8],c8,sum[8],c9);
full_adder fa10(x[9],y[9],c9,sum[9],c10);
full_adder fa11(x[10],y[10],c10,sum[10],c11);
full_adder fa12(x[11],y[11],c11,sum[11],c12);
full_adder fa13(x[12],y[12],c12,sum[12],c13);
full_adder fa14(x[13],y[13],c13,sum[13],c14);
full_adder fa15(x[14],y[14],c14,sum[14],c15);
full_adder fa16(x[15],y[15],c15,sum[15],c16);
full_adder fa17(x[16],y[16],c16,sum[16],c17);
full_adder fa18(x[17],y[17],c17,sum[17],c18);
full_adder fa19(x[18],y[18],c18,sum[18],c19);
full_adder fa20(x[19],y[19],c19,sum[19],c20);
full_adder fa21(x[20],y[20],c20,sum[20],c21);
full_adder fa22(x[21],y[21],c21,sum[21],c22);
full_adder fa23(x[22],y[22],c22,sum[22],c23);
full_adder fa24(x[23],y[23],c23,sum[23],c24);
full_adder fa25(x[24],y[24],c24,sum[24],c25);
full_adder fa26(x[25],y[25],c25,sum[25],c26);
full_adder fa27(x[26],y[26],c26,sum[26],c27);
full_adder fa28(x[27],y[27],c27,sum[27],c28);
full_adder fa29(x[28],y[28],c28,sum[28],c29);
full_adder fa30(x[29],y[29],c29,sum[29],c30);
full_adder fa31(x[30],y[30],c30,sum[30],c31);
full_adder fa32(x[31],y[31],c31,sum[31],ov);
xor(cout,c31,ov);
endmodule