module subop(difference, x, y,borrow);
input [31:0] x,y;
output borrow;
output [31:0] difference;
wire ov,c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29,c30,c31;

full_sub fs1(x[0],y[0],1'b0,difference[0],c1);
full_sub fs2(x[1],y[1],c1,difference[1],c2);
full_sub fs3(x[2],y[2],c2,difference[2],c3);
full_sub fs4(x[3],y[3],c3,difference[3],c4);
full_sub fs5(x[4],y[4],c4,difference[4],c5);
full_sub fs6(x[5],y[5],c5,difference[5],c6);
full_sub fs7(x[6],y[6],c6,difference[6],c7);
full_sub fs8(x[7],y[7],c7,difference[7],c8);
full_sub fs9(x[8],y[8],c8,difference[8],c9);
full_sub fs10(x[9],y[9],c9,difference[9],c10);
full_sub fs11(x[10],y[10],c10,difference[10],c11);
full_sub fs12(x[11],y[11],c11,difference[11],c12);
full_sub fs13(x[12],y[12],c12,difference[12],c13);
full_sub fs14(x[13],y[13],c13,difference[13],c14);
full_sub fs15(x[14],y[14],c14,difference[14],c15);
full_sub fs16(x[15],y[15],c15,difference[15],c16);
full_sub fs17(x[16],y[16],c16,difference[16],c17);
full_sub fs18(x[17],y[17],c17,difference[17],c18);
full_sub fs19(x[18],y[18],c18,difference[18],c19);
full_sub fs20(x[19],y[19],c19,difference[19],c20);
full_sub fs21(x[20],y[20],c20,difference[20],c21);
full_sub fs22(x[21],y[21],c21,difference[21],c22);
full_sub fs23(x[22],y[22],c22,difference[22],c23);
full_sub fs24(x[23],y[23],c23,difference[23],c24);
full_sub fs25(x[24],y[24],c24,difference[24],c25);
full_sub fs26(x[25],y[25],c25,difference[25],c26);
full_sub fs27(x[26],y[26],c26,difference[26],c27);
full_sub fs28(x[27],y[27],c27,difference[27],c28);
full_sub fs29(x[28],y[28],c28,difference[28],c29);
full_sub fs30(x[29],y[29],c29,difference[29],c30);
full_sub fs31(x[30],y[30],c30,difference[30],c31);
full_sub fs32(x[31],y[31],c31,difference[31],ov);
xor(borrow,c31,ov);
endmodule