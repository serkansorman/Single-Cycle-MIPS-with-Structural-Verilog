module shiftL(R, A, B, S);

input [31:0]  A;  
input [31:0]  B;
input S;  
output [31:0] R;

wire [31:0] s1,s2,s3,s4;


// 1 Bit Shift
mux2x1 m1(s1[0],A[0],S,B[0]);
mux2x1 m2(s1[1],A[1],A[0],B[0]);
mux2x1 m3(s1[2],A[2],A[1],B[0]);
mux2x1 m4(s1[3],A[3],A[2],B[0]);
mux2x1 m5(s1[4],A[4],A[3],B[0]);
mux2x1 m6(s1[5],A[5],A[4],B[0]);
mux2x1 m7(s1[6],A[6],A[5],B[0]);
mux2x1 m8(s1[7],A[7],A[6],B[0]);
mux2x1 m9(s1[8],A[8],A[7],B[0]);
mux2x1 m10(s1[9],A[9],A[8],B[0]);
mux2x1 m11(s1[10],A[10],A[9],B[0]);
mux2x1 m12(s1[11],A[11],A[10],B[0]);
mux2x1 m13(s1[12],A[12],A[11],B[0]);
mux2x1 m14(s1[13],A[13],A[12],B[0]);
mux2x1 m15(s1[14],A[14],A[13],B[0]);
mux2x1 m16(s1[15],A[15],A[14],B[0]);
mux2x1 m17(s1[16],A[16],A[15],B[0]);
mux2x1 m18(s1[17],A[17],A[16],B[0]);
mux2x1 m19(s1[18],A[18],A[17],B[0]);
mux2x1 m20(s1[19],A[19],A[18],B[0]);
mux2x1 m21(s1[20],A[20],A[19],B[0]);
mux2x1 m22(s1[21],A[21],A[20],B[0]);
mux2x1 m23(s1[22],A[22],A[21],B[0]);
mux2x1 m24(s1[23],A[23],A[22],B[0]);
mux2x1 m25(s1[24],A[24],A[23],B[0]);
mux2x1 m26(s1[25],A[25],A[24],B[0]);
mux2x1 m27(s1[26],A[26],A[25],B[0]);
mux2x1 m28(s1[27],A[27],A[26],B[0]);
mux2x1 m29(s1[28],A[28],A[27],B[0]);
mux2x1 m30(s1[29],A[29],A[28],B[0]);
mux2x1 m31(s1[30],A[30],A[29],B[0]);
mux2x1 m32(s1[31],A[31],A[30],B[0]);


//2 Bit Shift
mux2x1 m_1(s2[0],s1[0],S,B[1]);
mux2x1 m_2(s2[1],s1[1],S,B[1]);
mux2x1 m_3(s2[2],s1[2],s1[0],B[1]);
mux2x1 m_4(s2[3],s1[3],s1[1],B[1]);
mux2x1 m_5(s2[4],s1[4],s1[2],B[1]);
mux2x1 m_6(s2[5],s1[5],s1[3],B[1]);
mux2x1 m_7(s2[6],s1[6],s1[4],B[1]);
mux2x1 m_8(s2[7],s1[7],s1[5],B[1]);
mux2x1 m_9(s2[8],s1[8],s1[6],B[1]);
mux2x1 m_10(s2[9],s1[9],s1[7],B[1]);
mux2x1 m_11(s2[10],s1[10],s1[8],B[1]);
mux2x1 m_12(s2[11],s1[11],s1[9],B[1]);
mux2x1 m_13(s2[12],s1[12],s1[10],B[1]);
mux2x1 m_14(s2[13],s1[13],s1[11],B[1]);
mux2x1 m_15(s2[14],s1[14],s1[12],B[1]);
mux2x1 m_16(s2[15],s1[15],s1[13],B[1]);
mux2x1 m_17(s2[16],s1[16],s1[14],B[1]);
mux2x1 m_18(s2[17],s1[17],s1[15],B[1]);
mux2x1 m_19(s2[18],s1[18],s1[16],B[1]);
mux2x1 m_20(s2[19],s1[19],s1[17],B[1]);
mux2x1 m_21(s2[20],s1[20],s1[18],B[1]);
mux2x1 m_22(s2[21],s1[21],s1[19],B[1]);
mux2x1 m_23(s2[22],s1[22],s1[20],B[1]);
mux2x1 m_24(s2[23],s1[23],s1[21],B[1]);
mux2x1 m_25(s2[24],s1[24],s1[22],B[1]);
mux2x1 m_26(s2[25],s1[25],s1[23],B[1]);
mux2x1 m_27(s2[26],s1[26],s1[24],B[1]);
mux2x1 m_28(s2[27],s1[27],s1[25],B[1]);
mux2x1 m_29(s2[28],s1[28],s1[26],B[1]);
mux2x1 m_30(s2[29],s1[29],s1[27],B[1]);
mux2x1 m_31(s2[30],s1[30],s1[28],B[1]);
mux2x1 m_32(s2[31],s1[31],s1[29],B[1]);

//4 Bit Shift
mux2x1 m__1(s3[0],s2[0],S,B[2]);
mux2x1 m__2(s3[1],s2[1],S,B[2]);
mux2x1 m__3(s3[2],s2[2],S,B[2]);
mux2x1 m__4(s3[3],s2[3],S,B[2]);
mux2x1 m__5(s3[4],s2[4],s2[0],B[2]);
mux2x1 m__6(s3[5],s2[5],s2[1],B[2]);
mux2x1 m__7(s3[6],s2[6],s2[2],B[2]);
mux2x1 m__8(s3[7],s2[7],s2[3],B[2]);
mux2x1 m__9(s3[8],s2[8],s2[4],B[2]);
mux2x1 m__10(s3[9],s2[9],s2[5],B[2]);
mux2x1 m__11(s3[10],s2[10],s2[6],B[2]);
mux2x1 m__12(s3[11],s2[11],s2[7],B[2]);
mux2x1 m__13(s3[12],s2[12],s2[8],B[2]);
mux2x1 m__14(s3[13],s2[13],s2[9],B[2]);
mux2x1 m__15(s3[14],s2[14],s2[10],B[2]);
mux2x1 m__16(s3[15],s2[15],s2[11],B[2]);
mux2x1 m__17(s3[16],s2[16],s2[12],B[2]);
mux2x1 m__18(s3[17],s2[17],s2[13],B[2]);
mux2x1 m__19(s3[18],s2[18],s2[14],B[2]);
mux2x1 m__20(s3[19],s2[19],s2[15],B[2]);
mux2x1 m__21(s3[20],s2[20],s2[16],B[2]);
mux2x1 m__22(s3[21],s2[21],s2[17],B[2]);
mux2x1 m__23(s3[22],s2[22],s2[18],B[2]);
mux2x1 m__24(s3[23],s2[23],s2[19],B[2]);
mux2x1 m__25(s3[24],s2[24],s2[20],B[2]);
mux2x1 m__26(s3[25],s2[25],s2[21],B[2]);
mux2x1 m__27(s3[26],s2[26],s2[22],B[2]);
mux2x1 m__28(s3[27],s2[27],s2[23],B[2]);
mux2x1 m__29(s3[28],s2[28],s2[24],B[2]);
mux2x1 m__30(s3[29],s2[29],s2[25],B[2]);
mux2x1 m__31(s3[30],s2[30],s2[26],B[2]);
mux2x1 m__32(s3[31],s2[31],s2[27],B[2]);

//8 Bit Shift
mux2x1 m___1(s4[0],s3[0],S,B[3]);
mux2x1 m___2(s4[1],s3[1],S,B[3]);
mux2x1 m___3(s4[2],s3[2],S,B[3]);
mux2x1 m___4(s4[3],s3[3],S,B[3]);
mux2x1 m___5(s4[4],s3[4],S,B[3]);
mux2x1 m___6(s4[5],s3[5],S,B[3]);
mux2x1 m___7(s4[6],s3[6],S,B[3]);
mux2x1 m___8(s4[7],s3[7],S,B[3]);
mux2x1 m___9(s4[8],s3[8],s3[0],B[3]);
mux2x1 m___10(s4[9],s3[9],s3[1],B[3]);
mux2x1 m___11(s4[10],s3[10],s3[2],B[3]);
mux2x1 m___12(s4[11],s3[11],s3[3],B[3]);
mux2x1 m___13(s4[12],s3[12],s3[4],B[3]);
mux2x1 m___14(s4[13],s3[13],s3[5],B[3]);
mux2x1 m___15(s4[14],s3[14],s3[6],B[3]);
mux2x1 m___16(s4[15],s3[15],s3[7],B[3]);
mux2x1 m___17(s4[16],s3[16],s3[8],B[3]);
mux2x1 m___18(s4[17],s3[17],s3[9],B[3]);
mux2x1 m___19(s4[18],s3[18],s3[10],B[3]);
mux2x1 m___20(s4[19],s3[19],s3[11],B[3]);
mux2x1 m___21(s4[20],s3[20],s3[12],B[3]);
mux2x1 m___22(s4[21],s3[21],s3[13],B[3]);
mux2x1 m___23(s4[22],s3[22],s3[14],B[3]);
mux2x1 m___24(s4[23],s3[23],s3[15],B[3]);
mux2x1 m___25(s4[24],s3[24],s3[16],B[3]);
mux2x1 m___26(s4[25],s3[25],s3[17],B[3]);
mux2x1 m___27(s4[26],s3[26],s3[18],B[3]);
mux2x1 m___28(s4[27],s3[27],s3[19],B[3]);
mux2x1 m___29(s4[28],s3[28],s3[20],B[3]);
mux2x1 m___30(s4[29],s3[29],s3[21],B[3]);
mux2x1 m___31(s4[30],s3[30],s3[22],B[3]);
mux2x1 m___32(s4[31],s3[31],s3[23],B[3]);

//16 Bit Shift
mux2x1 m____1(R[0],s4[0],S,B[4]);
mux2x1 m____2(R[1],s4[1],S,B[4]);
mux2x1 m____3(R[2],s4[2],S,B[4]);
mux2x1 m____4(R[3],s4[3],S,B[4]);
mux2x1 m____5(R[4],s4[4],S,B[4]);
mux2x1 m____6(R[5],s4[5],S,B[4]);
mux2x1 m____7(R[6],s4[6],S,B[4]);
mux2x1 m____8(R[7],s4[7],S,B[4]);
mux2x1 m____9(R[8],s4[8],S,B[4]);
mux2x1 m____10(R[9],s4[9],S,B[4]);
mux2x1 m____11(R[10],s4[10],S,B[4]);
mux2x1 m____12(R[11],s4[11],S,B[4]);
mux2x1 m____13(R[12],s4[12],S,B[4]);
mux2x1 m____14(R[13],s4[13],S,B[4]);
mux2x1 m____15(R[14],s4[14],S,B[4]);
mux2x1 m____16(R[15],s4[15],S,B[4]);
mux2x1 m____17(R[16],s4[16],s4[0],B[4]);
mux2x1 m____18(R[17],s4[17],s4[1],B[4]);
mux2x1 m____19(R[18],s4[18],s4[2],B[4]);
mux2x1 m____20(R[19],s4[19],s4[3],B[4]);
mux2x1 m____21(R[20],s4[20],s4[4],B[4]);
mux2x1 m____22(R[21],s4[21],s4[5],B[4]);
mux2x1 m____23(R[22],s4[22],s4[6],B[4]);
mux2x1 m____24(R[23],s4[23],s4[7],B[4]);
mux2x1 m____25(R[24],s4[24],s4[8],B[4]);
mux2x1 m____26(R[25],s4[25],s4[9],B[4]);
mux2x1 m____27(R[26],s4[26],s4[10],B[4]);
mux2x1 m____28(R[27],s4[27],s4[11],B[4]);
mux2x1 m____29(R[28],s4[28],s4[12],B[4]);
mux2x1 m____30(R[29],s4[29],s4[13],B[4]);
mux2x1 m____31(R[30],s4[30],s4[14],B[4]);
mux2x1 m____32(R[31],s4[31],s4[15],B[4]);


endmodule