module mux8x1_32(out,a,b,c,d,e,f,g,h,s);
input [31:0] a,b,c,d,e,f,g,h;
input [2:0] s;
output[31:0] out;

mux8x1 mu1(out[0],a[0],b[0],c[0],d[0],e[0],f[0],g[0],h[0],s);
mux8x1 mu2(out[1],a[1],b[1],c[1],d[1],e[1],f[1],g[1],h[1],s);
mux8x1 mu3(out[2],a[2],b[2],c[2],d[2],e[2],f[2],g[2],h[2],s);
mux8x1 mu4(out[3],a[3],b[3],c[3],d[3],e[3],f[3],g[3],h[3],s);
mux8x1 mu5(out[4],a[4],b[4],c[4],d[4],e[4],f[4],g[4],h[4],s);
mux8x1 mu6(out[5],a[5],b[5],c[5],d[5],e[5],f[5],g[5],h[5],s);
mux8x1 mu7(out[6],a[6],b[6],c[6],d[6],e[6],f[6],g[6],h[6],s);
mux8x1 mu8(out[7],a[7],b[7],c[7],d[7],e[7],f[7],g[7],h[7],s);
mux8x1 mu9(out[8],a[8],b[8],c[8],d[8],e[8],f[8],g[8],h[8],s);
mux8x1 mu10(out[9],a[9],b[9],c[9],d[9],e[9],f[9],g[9],h[9],s);
mux8x1 mu11(out[10],a[10],b[10],c[10],d[10],e[10],f[10],g[10],h[10],s);
mux8x1 mu12(out[11],a[11],b[11],c[11],d[11],e[11],f[11],g[11],h[11],s);
mux8x1 mu13(out[12],a[12],b[12],c[12],d[12],e[12],f[12],g[12],h[12],s);
mux8x1 mu14(out[13],a[13],b[13],c[13],d[13],e[13],f[13],g[13],h[13],s);
mux8x1 mu15(out[14],a[14],b[14],c[14],d[14],e[14],f[14],g[14],h[14],s);
mux8x1 mu16(out[15],a[15],b[15],c[15],d[15],e[15],f[15],g[15],h[15],s);
mux8x1 mu17(out[16],a[16],b[16],c[16],d[16],e[16],f[16],g[16],h[16],s);
mux8x1 mu18(out[17],a[17],b[17],c[17],d[17],e[17],f[17],g[17],h[17],s);
mux8x1 mu19(out[18],a[18],b[18],c[18],d[18],e[18],f[18],g[18],h[18],s);
mux8x1 mu20(out[19],a[19],b[19],c[19],d[19],e[19],f[19],g[19],h[19],s);
mux8x1 mu21(out[20],a[20],b[20],c[20],d[20],e[20],f[20],g[20],h[20],s);
mux8x1 mu22(out[21],a[21],b[21],c[21],d[21],e[21],f[21],g[21],h[21],s);
mux8x1 mu23(out[22],a[22],b[22],c[22],d[22],e[22],f[22],g[22],h[22],s);
mux8x1 mu24(out[23],a[23],b[23],c[23],d[23],e[23],f[23],g[23],h[23],s);
mux8x1 mu25(out[24],a[24],b[24],c[24],d[24],e[24],f[24],g[24],h[24],s);
mux8x1 mu26(out[25],a[25],b[25],c[25],d[25],e[25],f[25],g[25],h[25],s);
mux8x1 mu27(out[26],a[26],b[26],c[26],d[26],e[26],f[26],g[26],h[26],s);
mux8x1 mu28(out[27],a[27],b[27],c[27],d[27],e[27],f[27],g[27],h[27],s);
mux8x1 mu29(out[28],a[28],b[28],c[28],d[28],e[28],f[28],g[28],h[28],s);
mux8x1 mu30(out[29],a[29],b[29],c[29],d[29],e[29],f[29],g[29],h[29],s);
mux8x1 mu31(out[30],a[30],b[30],c[30],d[30],e[30],f[30],g[30],h[30],s);
mux8x1 mu32(out[31],a[31],b[31],c[31],d[31],e[31],f[31],g[31],h[31],s);
endmodule