module mux2x1_32(out,a,b,s);
input [31:0] a,b;
input s;
output[31:0] out;

mux2x1 mu1(out[0],a[0],b[0],s);
mux2x1 mu2(out[1],a[1],b[1],s);
mux2x1 mu3(out[2],a[2],b[2],s);
mux2x1 mu4(out[3],a[3],b[3],s);
mux2x1 mu5(out[4],a[4],b[4],s);
mux2x1 mu6(out[5],a[5],b[5],s);
mux2x1 mu7(out[6],a[6],b[6],s);
mux2x1 mu8(out[7],a[7],b[7],s);
mux2x1 mu9(out[8],a[8],b[8],s);
mux2x1 mu10(out[9],a[9],b[9],s);
mux2x1 mu11(out[10],a[10],b[10],s);
mux2x1 mu12(out[11],a[11],b[11],s);
mux2x1 mu13(out[12],a[12],b[12],s);
mux2x1 mu14(out[13],a[13],b[13],s);
mux2x1 mu15(out[14],a[14],b[14],s);
mux2x1 mu16(out[15],a[15],b[15],s);
mux2x1 mu17(out[16],a[16],b[16],s);
mux2x1 mu18(out[17],a[17],b[17],s);
mux2x1 mu19(out[18],a[18],b[18],s);
mux2x1 mu20(out[19],a[19],b[19],s);
mux2x1 mu21(out[20],a[20],b[20],s);
mux2x1 mu22(out[21],a[21],b[21],s);
mux2x1 mu23(out[22],a[22],b[22],s);
mux2x1 mu24(out[23],a[23],b[23],s);
mux2x1 mu25(out[24],a[24],b[24],s);
mux2x1 mu26(out[25],a[25],b[25],s);
mux2x1 mu27(out[26],a[26],b[26],s);
mux2x1 mu28(out[27],a[27],b[27],s);
mux2x1 mu29(out[28],a[28],b[28],s);
mux2x1 mu30(out[29],a[29],b[29],s);
mux2x1 mu31(out[30],a[30],b[30],s);
mux2x1 mu32(out[31],a[31],b[31],s);
endmodule